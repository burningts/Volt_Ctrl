// nios.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module nios (
		input  wire        clk_clk,          //        clk.clk
		output wire        epcs_flash_dclk,  // epcs_flash.dclk
		output wire        epcs_flash_sce,   //           .sce
		output wire        epcs_flash_sdo,   //           .sdo
		input  wire        epcs_flash_data0, //           .data0
		output wire        ldac_n_export,    //     ldac_n.export
		output wire [31:0] oe_export,        //         oe.export
		output wire        pio_led_export,   //    pio_led.export
		input  wire        reset_reset_n,    //      reset.reset_n
		input  wire        spi_MISO,         //        spi.MISO
		output wire        spi_MOSI,         //           .MOSI
		output wire        spi_SCLK,         //           .SCLK
		output wire        spi_SS_n,         //           .SS_n
		input  wire        uart_rxd,         //       uart.rxd
		output wire        uart_txd          //           .txd
	);

	wire  [31:0] nios_data_master_readdata;                                 // mm_interconnect_0:nios_data_master_readdata -> nios:d_readdata
	wire         nios_data_master_waitrequest;                              // mm_interconnect_0:nios_data_master_waitrequest -> nios:d_waitrequest
	wire         nios_data_master_debugaccess;                              // nios:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios_data_master_debugaccess
	wire  [16:0] nios_data_master_address;                                  // nios:d_address -> mm_interconnect_0:nios_data_master_address
	wire   [3:0] nios_data_master_byteenable;                               // nios:d_byteenable -> mm_interconnect_0:nios_data_master_byteenable
	wire         nios_data_master_read;                                     // nios:d_read -> mm_interconnect_0:nios_data_master_read
	wire         nios_data_master_readdatavalid;                            // mm_interconnect_0:nios_data_master_readdatavalid -> nios:d_readdatavalid
	wire         nios_data_master_write;                                    // nios:d_write -> mm_interconnect_0:nios_data_master_write
	wire  [31:0] nios_data_master_writedata;                                // nios:d_writedata -> mm_interconnect_0:nios_data_master_writedata
	wire  [31:0] nios_instruction_master_readdata;                          // mm_interconnect_0:nios_instruction_master_readdata -> nios:i_readdata
	wire         nios_instruction_master_waitrequest;                       // mm_interconnect_0:nios_instruction_master_waitrequest -> nios:i_waitrequest
	wire  [16:0] nios_instruction_master_address;                           // nios:i_address -> mm_interconnect_0:nios_instruction_master_address
	wire         nios_instruction_master_read;                              // nios:i_read -> mm_interconnect_0:nios_instruction_master_read
	wire         nios_instruction_master_readdatavalid;                     // mm_interconnect_0:nios_instruction_master_readdatavalid -> nios:i_readdatavalid
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;       // mm_interconnect_0:jtag_avalon_jtag_slave_chipselect -> jtag:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;         // jtag:av_readdata -> mm_interconnect_0:jtag_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest;      // jtag:av_waitrequest -> mm_interconnect_0:jtag_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;          // mm_interconnect_0:jtag_avalon_jtag_slave_address -> jtag:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;             // mm_interconnect_0:jtag_avalon_jtag_slave_read -> jtag:av_read_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;            // mm_interconnect_0:jtag_avalon_jtag_slave_write -> jtag:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;        // mm_interconnect_0:jtag_avalon_jtag_slave_writedata -> jtag:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;            // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;             // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_nios_debug_mem_slave_readdata;           // nios:debug_mem_slave_readdata -> mm_interconnect_0:nios_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios_debug_mem_slave_waitrequest;        // nios:debug_mem_slave_waitrequest -> mm_interconnect_0:nios_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios_debug_mem_slave_debugaccess;        // mm_interconnect_0:nios_debug_mem_slave_debugaccess -> nios:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios_debug_mem_slave_address;            // mm_interconnect_0:nios_debug_mem_slave_address -> nios:debug_mem_slave_address
	wire         mm_interconnect_0_nios_debug_mem_slave_read;               // mm_interconnect_0:nios_debug_mem_slave_read -> nios:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios_debug_mem_slave_byteenable;         // mm_interconnect_0:nios_debug_mem_slave_byteenable -> nios:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios_debug_mem_slave_write;              // mm_interconnect_0:nios_debug_mem_slave_write -> nios:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios_debug_mem_slave_writedata;          // mm_interconnect_0:nios_debug_mem_slave_writedata -> nios:debug_mem_slave_writedata
	wire         mm_interconnect_0_epcs_flash_epcs_control_port_chipselect; // mm_interconnect_0:epcs_flash_epcs_control_port_chipselect -> epcs_flash:chipselect
	wire  [31:0] mm_interconnect_0_epcs_flash_epcs_control_port_readdata;   // epcs_flash:readdata -> mm_interconnect_0:epcs_flash_epcs_control_port_readdata
	wire   [8:0] mm_interconnect_0_epcs_flash_epcs_control_port_address;    // mm_interconnect_0:epcs_flash_epcs_control_port_address -> epcs_flash:address
	wire         mm_interconnect_0_epcs_flash_epcs_control_port_read;       // mm_interconnect_0:epcs_flash_epcs_control_port_read -> epcs_flash:read_n
	wire         mm_interconnect_0_epcs_flash_epcs_control_port_write;      // mm_interconnect_0:epcs_flash_epcs_control_port_write -> epcs_flash:write_n
	wire  [31:0] mm_interconnect_0_epcs_flash_epcs_control_port_writedata;  // mm_interconnect_0:epcs_flash_epcs_control_port_writedata -> epcs_flash:writedata
	wire         mm_interconnect_0_rom_s1_chipselect;                       // mm_interconnect_0:rom_s1_chipselect -> rom:chipselect
	wire  [31:0] mm_interconnect_0_rom_s1_readdata;                         // rom:readdata -> mm_interconnect_0:rom_s1_readdata
	wire         mm_interconnect_0_rom_s1_debugaccess;                      // mm_interconnect_0:rom_s1_debugaccess -> rom:debugaccess
	wire  [11:0] mm_interconnect_0_rom_s1_address;                          // mm_interconnect_0:rom_s1_address -> rom:address
	wire   [3:0] mm_interconnect_0_rom_s1_byteenable;                       // mm_interconnect_0:rom_s1_byteenable -> rom:byteenable
	wire         mm_interconnect_0_rom_s1_write;                            // mm_interconnect_0:rom_s1_write -> rom:write
	wire  [31:0] mm_interconnect_0_rom_s1_writedata;                        // mm_interconnect_0:rom_s1_writedata -> rom:writedata
	wire         mm_interconnect_0_rom_s1_clken;                            // mm_interconnect_0:rom_s1_clken -> rom:clken
	wire         mm_interconnect_0_ram_s1_chipselect;                       // mm_interconnect_0:ram_s1_chipselect -> ram:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                         // ram:readdata -> mm_interconnect_0:ram_s1_readdata
	wire  [11:0] mm_interconnect_0_ram_s1_address;                          // mm_interconnect_0:ram_s1_address -> ram:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                       // mm_interconnect_0:ram_s1_byteenable -> ram:byteenable
	wire         mm_interconnect_0_ram_s1_write;                            // mm_interconnect_0:ram_s1_write -> ram:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                        // mm_interconnect_0:ram_s1_writedata -> ram:writedata
	wire         mm_interconnect_0_ram_s1_clken;                            // mm_interconnect_0:ram_s1_clken -> ram:clken
	wire         mm_interconnect_0_pio_oe_s1_chipselect;                    // mm_interconnect_0:pio_oe_s1_chipselect -> pio_oe:chipselect
	wire  [31:0] mm_interconnect_0_pio_oe_s1_readdata;                      // pio_oe:readdata -> mm_interconnect_0:pio_oe_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_oe_s1_address;                       // mm_interconnect_0:pio_oe_s1_address -> pio_oe:address
	wire         mm_interconnect_0_pio_oe_s1_write;                         // mm_interconnect_0:pio_oe_s1_write -> pio_oe:write_n
	wire  [31:0] mm_interconnect_0_pio_oe_s1_writedata;                     // mm_interconnect_0:pio_oe_s1_writedata -> pio_oe:writedata
	wire         mm_interconnect_0_pio_ldac_n_s1_chipselect;                // mm_interconnect_0:pio_ldac_n_s1_chipselect -> pio_ldac_n:chipselect
	wire  [31:0] mm_interconnect_0_pio_ldac_n_s1_readdata;                  // pio_ldac_n:readdata -> mm_interconnect_0:pio_ldac_n_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_ldac_n_s1_address;                   // mm_interconnect_0:pio_ldac_n_s1_address -> pio_ldac_n:address
	wire         mm_interconnect_0_pio_ldac_n_s1_write;                     // mm_interconnect_0:pio_ldac_n_s1_write -> pio_ldac_n:write_n
	wire  [31:0] mm_interconnect_0_pio_ldac_n_s1_writedata;                 // mm_interconnect_0:pio_ldac_n_s1_writedata -> pio_ldac_n:writedata
	wire         mm_interconnect_0_uart_s1_chipselect;                      // mm_interconnect_0:uart_s1_chipselect -> uart:chipselect
	wire  [15:0] mm_interconnect_0_uart_s1_readdata;                        // uart:readdata -> mm_interconnect_0:uart_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_s1_address;                         // mm_interconnect_0:uart_s1_address -> uart:address
	wire         mm_interconnect_0_uart_s1_read;                            // mm_interconnect_0:uart_s1_read -> uart:read_n
	wire         mm_interconnect_0_uart_s1_begintransfer;                   // mm_interconnect_0:uart_s1_begintransfer -> uart:begintransfer
	wire         mm_interconnect_0_uart_s1_write;                           // mm_interconnect_0:uart_s1_write -> uart:write_n
	wire  [15:0] mm_interconnect_0_uart_s1_writedata;                       // mm_interconnect_0:uart_s1_writedata -> uart:writedata
	wire         mm_interconnect_0_pio_led_s1_chipselect;                   // mm_interconnect_0:pio_led_s1_chipselect -> pio_led:chipselect
	wire  [31:0] mm_interconnect_0_pio_led_s1_readdata;                     // pio_led:readdata -> mm_interconnect_0:pio_led_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_led_s1_address;                      // mm_interconnect_0:pio_led_s1_address -> pio_led:address
	wire         mm_interconnect_0_pio_led_s1_write;                        // mm_interconnect_0:pio_led_s1_write -> pio_led:write_n
	wire  [31:0] mm_interconnect_0_pio_led_s1_writedata;                    // mm_interconnect_0:pio_led_s1_writedata -> pio_led:writedata
	wire         mm_interconnect_0_spi_spi_control_port_chipselect;         // mm_interconnect_0:spi_spi_control_port_chipselect -> spi:spi_select
	wire  [15:0] mm_interconnect_0_spi_spi_control_port_readdata;           // spi:data_to_cpu -> mm_interconnect_0:spi_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_spi_spi_control_port_address;            // mm_interconnect_0:spi_spi_control_port_address -> spi:mem_addr
	wire         mm_interconnect_0_spi_spi_control_port_read;               // mm_interconnect_0:spi_spi_control_port_read -> spi:read_n
	wire         mm_interconnect_0_spi_spi_control_port_write;              // mm_interconnect_0:spi_spi_control_port_write -> spi:write_n
	wire  [15:0] mm_interconnect_0_spi_spi_control_port_writedata;          // mm_interconnect_0:spi_spi_control_port_writedata -> spi:data_from_cpu
	wire         irq_mapper_receiver0_irq;                                  // jtag:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // spi:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                  // uart:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                  // epcs_flash:irq -> irq_mapper:receiver3_irq
	wire  [31:0] nios_irq_irq;                                              // irq_mapper:sender_irq -> nios:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [epcs_flash:reset_n, irq_mapper:reset, jtag:rst_n, mm_interconnect_0:nios_reset_reset_bridge_in_reset_reset, nios:reset_n, pio_ldac_n:reset_n, pio_led:reset_n, pio_oe:reset_n, ram:reset, rom:reset, rst_translator:in_reset, spi:reset_n, sysid:reset_n, uart:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [epcs_flash:reset_req, nios:reset_req, ram:reset_req, rom:reset_req, rst_translator:reset_req_in]
	wire         nios_debug_reset_request_reset;                            // nios:debug_reset_request -> rst_controller:reset_in1

	nios_epcs_flash epcs_flash (
		.clk        (clk_clk),                                                   //               clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.reset_req  (rst_controller_reset_out_reset_req),                        //                  .reset_req
		.address    (mm_interconnect_0_epcs_flash_epcs_control_port_address),    // epcs_control_port.address
		.chipselect (mm_interconnect_0_epcs_flash_epcs_control_port_chipselect), //                  .chipselect
		.read_n     (~mm_interconnect_0_epcs_flash_epcs_control_port_read),      //                  .read_n
		.readdata   (mm_interconnect_0_epcs_flash_epcs_control_port_readdata),   //                  .readdata
		.write_n    (~mm_interconnect_0_epcs_flash_epcs_control_port_write),     //                  .write_n
		.writedata  (mm_interconnect_0_epcs_flash_epcs_control_port_writedata),  //                  .writedata
		.irq        (irq_mapper_receiver3_irq),                                  //               irq.irq
		.dclk       (epcs_flash_dclk),                                           //          external.export
		.sce        (epcs_flash_sce),                                            //                  .export
		.sdo        (epcs_flash_sdo),                                            //                  .export
		.data0      (epcs_flash_data0)                                           //                  .export
	);

	nios_jtag jtag (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                              //               irq.irq
	);

	nios_nios nios (
		.clk                                 (clk_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                    //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                 //                          .reset_req
		.d_address                           (nios_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios_data_master_read),                              //                          .read
		.d_readdata                          (nios_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios_data_master_write),                             //                          .write
		.d_writedata                         (nios_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios_instruction_master_read),                       //                          .read
		.i_readdata                          (nios_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                    // custom_instruction_master.readra
	);

	nios_pio_ldac_n pio_ldac_n (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_pio_ldac_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_ldac_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_ldac_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_ldac_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_ldac_n_s1_readdata),   //                    .readdata
		.out_port   (ldac_n_export)                               // external_connection.export
	);

	nios_pio_ldac_n pio_led (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_pio_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_led_s1_readdata),   //                    .readdata
		.out_port   (pio_led_export)                           // external_connection.export
	);

	nios_pio_oe pio_oe (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_pio_oe_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_oe_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_oe_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_oe_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_oe_s1_readdata),   //                    .readdata
		.out_port   (oe_export)                               // external_connection.export
	);

	nios_ram ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	nios_rom rom (
		.clk         (clk_clk),                              //   clk1.clk
		.address     (mm_interconnect_0_rom_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_rom_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_rom_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_rom_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_rom_s1_write),       //       .write
		.readdata    (mm_interconnect_0_rom_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_rom_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_rom_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),       // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),   //       .reset_req
		.freeze      (1'b0)                                  // (terminated)
	);

	nios_spi spi (
		.clk           (clk_clk),                                           //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                   //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_spi_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_spi_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_spi_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_spi_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_spi_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_spi_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver1_irq),                          //              irq.irq
		.MISO          (spi_MISO),                                          //         external.export
		.MOSI          (spi_MOSI),                                          //                 .export
		.SCLK          (spi_SCLK),                                          //                 .export
		.SS_n          (spi_SS_n)                                           //                 .export
	);

	nios_sysid sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	nios_uart uart (
		.clk           (clk_clk),                                 //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address       (mm_interconnect_0_uart_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_s1_readdata),      //                    .readdata
		.rxd           (uart_rxd),                                // external_connection.export
		.txd           (uart_txd),                                //                    .export
		.irq           (irq_mapper_receiver2_irq)                 //                 irq.irq
	);

	nios_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                           (clk_clk),                                                   //                        clk_0_clk.clk
		.nios_reset_reset_bridge_in_reset_reset  (rst_controller_reset_out_reset),                            // nios_reset_reset_bridge_in_reset.reset
		.nios_data_master_address                (nios_data_master_address),                                  //                 nios_data_master.address
		.nios_data_master_waitrequest            (nios_data_master_waitrequest),                              //                                 .waitrequest
		.nios_data_master_byteenable             (nios_data_master_byteenable),                               //                                 .byteenable
		.nios_data_master_read                   (nios_data_master_read),                                     //                                 .read
		.nios_data_master_readdata               (nios_data_master_readdata),                                 //                                 .readdata
		.nios_data_master_readdatavalid          (nios_data_master_readdatavalid),                            //                                 .readdatavalid
		.nios_data_master_write                  (nios_data_master_write),                                    //                                 .write
		.nios_data_master_writedata              (nios_data_master_writedata),                                //                                 .writedata
		.nios_data_master_debugaccess            (nios_data_master_debugaccess),                              //                                 .debugaccess
		.nios_instruction_master_address         (nios_instruction_master_address),                           //          nios_instruction_master.address
		.nios_instruction_master_waitrequest     (nios_instruction_master_waitrequest),                       //                                 .waitrequest
		.nios_instruction_master_read            (nios_instruction_master_read),                              //                                 .read
		.nios_instruction_master_readdata        (nios_instruction_master_readdata),                          //                                 .readdata
		.nios_instruction_master_readdatavalid   (nios_instruction_master_readdatavalid),                     //                                 .readdatavalid
		.epcs_flash_epcs_control_port_address    (mm_interconnect_0_epcs_flash_epcs_control_port_address),    //     epcs_flash_epcs_control_port.address
		.epcs_flash_epcs_control_port_write      (mm_interconnect_0_epcs_flash_epcs_control_port_write),      //                                 .write
		.epcs_flash_epcs_control_port_read       (mm_interconnect_0_epcs_flash_epcs_control_port_read),       //                                 .read
		.epcs_flash_epcs_control_port_readdata   (mm_interconnect_0_epcs_flash_epcs_control_port_readdata),   //                                 .readdata
		.epcs_flash_epcs_control_port_writedata  (mm_interconnect_0_epcs_flash_epcs_control_port_writedata),  //                                 .writedata
		.epcs_flash_epcs_control_port_chipselect (mm_interconnect_0_epcs_flash_epcs_control_port_chipselect), //                                 .chipselect
		.jtag_avalon_jtag_slave_address          (mm_interconnect_0_jtag_avalon_jtag_slave_address),          //           jtag_avalon_jtag_slave.address
		.jtag_avalon_jtag_slave_write            (mm_interconnect_0_jtag_avalon_jtag_slave_write),            //                                 .write
		.jtag_avalon_jtag_slave_read             (mm_interconnect_0_jtag_avalon_jtag_slave_read),             //                                 .read
		.jtag_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),         //                                 .readdata
		.jtag_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),        //                                 .writedata
		.jtag_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest),      //                                 .waitrequest
		.jtag_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),       //                                 .chipselect
		.nios_debug_mem_slave_address            (mm_interconnect_0_nios_debug_mem_slave_address),            //             nios_debug_mem_slave.address
		.nios_debug_mem_slave_write              (mm_interconnect_0_nios_debug_mem_slave_write),              //                                 .write
		.nios_debug_mem_slave_read               (mm_interconnect_0_nios_debug_mem_slave_read),               //                                 .read
		.nios_debug_mem_slave_readdata           (mm_interconnect_0_nios_debug_mem_slave_readdata),           //                                 .readdata
		.nios_debug_mem_slave_writedata          (mm_interconnect_0_nios_debug_mem_slave_writedata),          //                                 .writedata
		.nios_debug_mem_slave_byteenable         (mm_interconnect_0_nios_debug_mem_slave_byteenable),         //                                 .byteenable
		.nios_debug_mem_slave_waitrequest        (mm_interconnect_0_nios_debug_mem_slave_waitrequest),        //                                 .waitrequest
		.nios_debug_mem_slave_debugaccess        (mm_interconnect_0_nios_debug_mem_slave_debugaccess),        //                                 .debugaccess
		.pio_ldac_n_s1_address                   (mm_interconnect_0_pio_ldac_n_s1_address),                   //                    pio_ldac_n_s1.address
		.pio_ldac_n_s1_write                     (mm_interconnect_0_pio_ldac_n_s1_write),                     //                                 .write
		.pio_ldac_n_s1_readdata                  (mm_interconnect_0_pio_ldac_n_s1_readdata),                  //                                 .readdata
		.pio_ldac_n_s1_writedata                 (mm_interconnect_0_pio_ldac_n_s1_writedata),                 //                                 .writedata
		.pio_ldac_n_s1_chipselect                (mm_interconnect_0_pio_ldac_n_s1_chipselect),                //                                 .chipselect
		.pio_led_s1_address                      (mm_interconnect_0_pio_led_s1_address),                      //                       pio_led_s1.address
		.pio_led_s1_write                        (mm_interconnect_0_pio_led_s1_write),                        //                                 .write
		.pio_led_s1_readdata                     (mm_interconnect_0_pio_led_s1_readdata),                     //                                 .readdata
		.pio_led_s1_writedata                    (mm_interconnect_0_pio_led_s1_writedata),                    //                                 .writedata
		.pio_led_s1_chipselect                   (mm_interconnect_0_pio_led_s1_chipselect),                   //                                 .chipselect
		.pio_oe_s1_address                       (mm_interconnect_0_pio_oe_s1_address),                       //                        pio_oe_s1.address
		.pio_oe_s1_write                         (mm_interconnect_0_pio_oe_s1_write),                         //                                 .write
		.pio_oe_s1_readdata                      (mm_interconnect_0_pio_oe_s1_readdata),                      //                                 .readdata
		.pio_oe_s1_writedata                     (mm_interconnect_0_pio_oe_s1_writedata),                     //                                 .writedata
		.pio_oe_s1_chipselect                    (mm_interconnect_0_pio_oe_s1_chipselect),                    //                                 .chipselect
		.ram_s1_address                          (mm_interconnect_0_ram_s1_address),                          //                           ram_s1.address
		.ram_s1_write                            (mm_interconnect_0_ram_s1_write),                            //                                 .write
		.ram_s1_readdata                         (mm_interconnect_0_ram_s1_readdata),                         //                                 .readdata
		.ram_s1_writedata                        (mm_interconnect_0_ram_s1_writedata),                        //                                 .writedata
		.ram_s1_byteenable                       (mm_interconnect_0_ram_s1_byteenable),                       //                                 .byteenable
		.ram_s1_chipselect                       (mm_interconnect_0_ram_s1_chipselect),                       //                                 .chipselect
		.ram_s1_clken                            (mm_interconnect_0_ram_s1_clken),                            //                                 .clken
		.rom_s1_address                          (mm_interconnect_0_rom_s1_address),                          //                           rom_s1.address
		.rom_s1_write                            (mm_interconnect_0_rom_s1_write),                            //                                 .write
		.rom_s1_readdata                         (mm_interconnect_0_rom_s1_readdata),                         //                                 .readdata
		.rom_s1_writedata                        (mm_interconnect_0_rom_s1_writedata),                        //                                 .writedata
		.rom_s1_byteenable                       (mm_interconnect_0_rom_s1_byteenable),                       //                                 .byteenable
		.rom_s1_chipselect                       (mm_interconnect_0_rom_s1_chipselect),                       //                                 .chipselect
		.rom_s1_clken                            (mm_interconnect_0_rom_s1_clken),                            //                                 .clken
		.rom_s1_debugaccess                      (mm_interconnect_0_rom_s1_debugaccess),                      //                                 .debugaccess
		.spi_spi_control_port_address            (mm_interconnect_0_spi_spi_control_port_address),            //             spi_spi_control_port.address
		.spi_spi_control_port_write              (mm_interconnect_0_spi_spi_control_port_write),              //                                 .write
		.spi_spi_control_port_read               (mm_interconnect_0_spi_spi_control_port_read),               //                                 .read
		.spi_spi_control_port_readdata           (mm_interconnect_0_spi_spi_control_port_readdata),           //                                 .readdata
		.spi_spi_control_port_writedata          (mm_interconnect_0_spi_spi_control_port_writedata),          //                                 .writedata
		.spi_spi_control_port_chipselect         (mm_interconnect_0_spi_spi_control_port_chipselect),         //                                 .chipselect
		.sysid_control_slave_address             (mm_interconnect_0_sysid_control_slave_address),             //              sysid_control_slave.address
		.sysid_control_slave_readdata            (mm_interconnect_0_sysid_control_slave_readdata),            //                                 .readdata
		.uart_s1_address                         (mm_interconnect_0_uart_s1_address),                         //                          uart_s1.address
		.uart_s1_write                           (mm_interconnect_0_uart_s1_write),                           //                                 .write
		.uart_s1_read                            (mm_interconnect_0_uart_s1_read),                            //                                 .read
		.uart_s1_readdata                        (mm_interconnect_0_uart_s1_readdata),                        //                                 .readdata
		.uart_s1_writedata                       (mm_interconnect_0_uart_s1_writedata),                       //                                 .writedata
		.uart_s1_begintransfer                   (mm_interconnect_0_uart_s1_begintransfer),                   //                                 .begintransfer
		.uart_s1_chipselect                      (mm_interconnect_0_uart_s1_chipselect)                       //                                 .chipselect
	);

	nios_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (nios_irq_irq)                    //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios_debug_reset_request_reset),     // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
